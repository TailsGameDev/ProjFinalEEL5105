library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity decod_nv is
port (
		G: in std_logic_vector(1 downto 0);
		D: out std_logic_vector(6 downto 0);
		enable: in std_logic
       );
end decod_nv;

architecture circuito of decod_nv is
begin
	D <=	"1111111" when enable = '0' else
			"1111001" when G = "00" else
			"0100100" when G = "01" else
			"0110000" when G = "10" else
			"0011001" when G = "11" else
			"1111111";
end circuito;